/*#####################################################################################################################################
## Package name : project_pkg
## Revision     : 
## Release note :   
/*#####################################################################################################################################*/

package project_pkg ;

  typedef class Transaction ;
  typedef class Driver;
  typedef class Sequencer;

  `include "transaction.svh"
  `include "driver.svh"
  `include "sequencer.svh"




endpackage