/*#####################################################################################################################################
## Package name : project_pkg
## Revision     : 
## Release note :   
/*#####################################################################################################################################*/

package project_pkg ;

  typedef class Transaction ;
  typedef class Driver;
  `include "transaction.svh"
  `include "driver.svh"




endpackage