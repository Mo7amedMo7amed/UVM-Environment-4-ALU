module alu (
	input rst_n, alu_clk, alu_enable_a, alu_enable_b, alu_enable, alu_irq_clr,
	input [7:0] alu_in_a, alu_in_b,
	input [1:0] alu_op_a, alu_op_b,
	output [7:0] alu_out,
	output alu_irq
);





endmodule