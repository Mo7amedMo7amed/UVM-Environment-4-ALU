package project_pkg ;
typedef class Transaction ;
`include "transaction.svh"




endpackage