/*#####################################################################################################################################
## Class name     : Monitor
## Revision       : 
## Release note   :   
/*#####################################################################################################################################*/

import uvm_pkg::*;
`include "uvm_macros.svh"
import project_pkg::*;

`ifndef Monitor_exists
`define Monitor_exists
class Monitor extends uvm_monitor ;





endclass
`endif 